* Circuit: Empty Circuit


.end