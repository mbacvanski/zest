.title NewAPICircuit

V1 vin gnd DC 12.0
R1 vin vout 10000.0
R2 vout n1 5000.0

.end