* Circuit: MultiInstanceTest

* ===== Subcircuit Definitions ===== *
.SUBCKT VOLTAGE_DIVIDER vin vout gnd
R1 vin vout 10000
R2 vout gnd 10000
.ENDS VOLTAGE_DIVIDER

* ===== Main Circuit Components ===== *
V1 N1 N2 DC 15.0
XU1 N1 N3 N2 VOLTAGE_DIVIDER
XU2 N3 N4 N2 VOLTAGE_DIVIDER

.end