* Circuit: Voltage Divider

V1 N1 gnd DC 12.0
R1 N1 N2 1000
R2 N2 gnd 2000

.end