* Circuit: Netlist Test

V1 V1_pos gnd DC 15.0
R1 V1_pos R1_n2 1500
R2 R1_n2 gnd 3000

.end