* Circuit: RC Filter

V1 R1_n1 gnd DC 5.0
R1 R1_n1 C1_pos 1000
C1 C1_pos gnd 1e-06

.end