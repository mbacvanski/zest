* Circuit: Mixed_Subcircuit_Types_Test

* ===== Model Includes ===== *
.INCLUDE "/Users/marc/Code/zest/tests/models/custom_resistor.lib"

* ===== Subcircuit Definitions ===== *
.SUBCKT RC_FILTER_STAGE_CUSTOM vin vout gnd
XR_custom vin vout CUSTOM_RESISTOR
CC_internal vout gnd 1e-06
.ENDS RC_FILTER_STAGE_CUSTOM

.SUBCKT VOLTAGE_DIVIDER_CUSTOM vin vout gnd
XR1_custom vin vout CUSTOM_RESISTOR
XR2_custom vout gnd CUSTOM_RESISTOR
.ENDS VOLTAGE_DIVIDER_CUSTOM

* ===== Main Circuit Components ===== *
V1 N1 gnd DC 5.0
XX_RC_Filter N1 N2 gnd RC_FILTER_STAGE_CUSTOM
XX_Voltage_Divider N2 N3 gnd VOLTAGE_DIVIDER_CUSTOM

* Initial Conditions
.IC V(N2)=0.0
.IC V(N3)=0.0

.end