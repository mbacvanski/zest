* Circuit: Simple Circuit

V1 R1_n1 gnd DC 5.0
R1 R1_n1 gnd 1000

.end