* Circuit: Netlist Test

V1 N1 gnd DC 15.0
R1 N1 N2 1500
R2 N2 gnd 3000

.end