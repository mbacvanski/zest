* Circuit: Simple Circuit

V1 V1_pos gnd DC 5.0
R1 V1_pos gnd 1000

.end