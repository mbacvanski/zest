* Circuit: Disconnected Test

V1 N1 N2 DC 5.0
R1 N3 N4 1000

.end