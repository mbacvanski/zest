* Circuit: Simple Circuit

V1 N1 gnd DC 5.0
R1 N1 gnd 1000

.end