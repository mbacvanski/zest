* Circuit: Voltage Divider

V1 V1_pos gnd DC 12.0
R1 V1_pos R1_n2 1000
R2 R1_n2 gnd 2000

.end