* Circuit: RC Filter

V1 N1 gnd DC 5.0
R1 N1 N2 1000
C1 N2 gnd 1e-06

.end